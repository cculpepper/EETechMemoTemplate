** Profile: "SCHEMATIC1-bnjkj"  [ C:\USERS\FPS7806\DESKTOP\lab02\lab2-PSpiceFiles\SCHEMATIC1\bnjkj.sim ] 

** Creating circuit file "bnjkj.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../lab2-pspicefiles/lab2.lib" 
* From [PSPICE NETLIST] section of C:\Users\fps7806\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 
.STEP LIN PARAM RVAL 1000 2500 500 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
